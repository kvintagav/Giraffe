module control_reg(
input wire CLK,
input wire [`FSMC_WIDTH-1:0] START_ADDR,
input wire [`FSMC_WIDTH-1:0] MOUNT_BYTE,
input wire READ,
input wire WRITE


);

endmodule
